'''***\$._svg_xmlv-version="1.1"/encoding="utf-8"/>
# Generator: Adobe Illustrator 16.0.0, SVG Export Plug-In . SVG Version: 6.00 Build #2)  -->
'DOCTYPE svg PUBLIC "-//W3C//DTD SVG 1.1//EN" "http://www.w3.org/Graphics/SVG/1.1/DTD/svg11.dtd">
<svg version="1.1" id="Layer_1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
	 width="2321.52px" height="432.99px" viewBox="0 0 2321.52 432.99" enable-background="new 0 0 2321.52 432.99"
	 xml:space="preserve">
<g>
	<g>
		<g>
			<path fill="#FC7E00" d="M198.143,355.152l7.171-15.141l11.02,5.204l2.822-5.988l-9.407-12.745l-16.688-7.908l-6.046,12.766
				l11.016,5.222l-8.804,18.591h-5.153c-2.334-5.252-2.442-6.829-3.365-8.112c-1.034-1.441-2.771-2.028-4.135-1.496l-2.538-3.527
				l2.022-1.463l-4.332-6.045l-4.061,2.9l-8.298-11.578l-3.545-8.298l-5.394-3.661l-3.67,2.63l1.747,6.286l6.724,6.018l8.301,11.575
				l-4.047,2.907l4.35,6.046l2.021-1.452l2.531,3.531c-0.804,0.967-0.879,2.426-0.245,3.739h-27.927v-8.601
				c4.98-2.534,8.417-7.69,8.417-13.672c0-6.52-4.075-12.08-9.801-14.306v15.693h-11.08v-15.693
				c-5.733,2.226-9.797,7.786-9.797,14.306c0,5.981,3.426,11.138,8.41,13.672v8.601h-18.343v22.396h121.077v-22.396H198.143z"/>
			<rect x="108.018" y="383.163" fill="#FC7E00" width="121.077" height="44.689"/>
		</g>
		<path fill="#FC7E00" d="M261.856,5.137H75.26c-37.86,0-68.551,30.691-68.551,68.559v285.615c0,37.85,30.691,68.541,68.551,68.541
			h4.953h9.686h4.163v-72.7h-4.176h-9.672H59.879V77.841H277.23v277.311h-17.535h-10.673h-5.971v72.7h5.957h10.687h2.161
			c37.856,0,68.548-30.691,68.548-68.541V73.696C330.404,35.829,299.713,5.137,261.856,5.137z"/>
	</g>
	<g>
		<path fill="#FC7E00" d="M380.54,299.004V132.809h31.961l56.373,126.096l55.205-126.096h30.792v166.195h-28.473V183.247
			l-45.097,115.758h-26.264l-46.02-115.758v115.758H380.54z"/>
		<path fill="#FC7E00" d="M581.023,237.999c0-40.91,20.146-61.365,60.433-61.365c40.296,0,60.442,20.455,60.442,61.365
			c0,40.828-20.146,61.24-60.442,61.24C601.327,299.239,581.182,278.827,581.023,237.999z M641.456,275.772
			c19.76,0,29.64-12.75,29.64-38.244c0-24.877-9.88-37.304-29.64-37.304c-19.758,0-29.632,12.427-29.632,37.304
			C611.824,263.022,621.698,275.772,641.456,275.772z"/>
		<path fill="#FC7E00" d="M725.143,132.809h30.793v53.462c9.226-6.199,19.487-9.295,30.799-9.295
			c34.717,0,52.072,19.532,52.072,58.577c0,42.307-19.877,63.451-59.627,63.451c-16.731,0-34.75-1.658-54.037-4.99V132.809z
			 M755.936,270.77c7.05,2.242,15.228,3.371,24.523,3.371c18.596,0,27.892-13.135,27.892-39.4c0-21.466-8.018-32.197-24.054-32.197
			c-10.388,0-19.834,2.099-28.361,6.286V270.77z"/>
		<path fill="#FC7E00" d="M892.844,132.809v24.403h-30.791v-24.403H892.844z M892.844,176.976v122.028h-30.791V176.976H892.844z"/>
		<path fill="#FC7E00" d="M952.702,132.809v166.195h-30.798V132.809H952.702z"/>
		<path fill="#FC7E00" d="M1033.241,176.976c37.036,0,55.558,18.91,55.558,56.712c0,5.041-0.353,10.084-1.052,15.113h-81.004
			c0,17.209,12.629,25.795,37.893,25.795c12.319,0,24.638-1.16,36.952-3.477v24.406c-10.768,2.316-23.86,3.479-39.279,3.479
			c-44.241,0-66.368-20.803-66.368-62.404C975.94,196.854,995.043,176.976,1033.241,176.976z M1006.743,227.415h52.069v-0.918
			c0-16.895-8.521-25.35-25.571-25.35C1016.969,201.147,1008.136,209.904,1006.743,227.415z"/>
		<path fill="#FC7E00" d="M1167.121,299.004V132.809h77.873c31.615,0,47.43,12.897,47.43,38.711
			c0,18.897-10.306,32.417-30.926,40.553c22.002,4.117,33.012,16.699,33.012,37.775c0,32.773-17.32,49.156-51.946,49.156H1167.121z
			 M1241.277,272.28c13.634,0,20.455-6.975,20.455-20.928c0-17.275-10.192-25.91-30.563-25.91h-9.296v-19.873
			c25.565-4.271,38.343-14.96,38.343-32.071c0-9.31-5.721-13.949-17.182-13.949h-45.11V272.28H1241.277z"/>
		<path fill="#FC7E00" d="M1427.584,176.976v122.028h-24.061l-3.727-15.564c-14.006,10.387-28.895,15.564-44.613,15.564
			c-24.958,0-37.43-14.752-37.43-44.281v-77.747h30.799v76.948c0,13.475,5.885,20.217,17.665,20.217
			c9.988,0,20.181-3.988,30.567-11.973v-85.192H1427.584z"/>
		<path fill="#FC7E00" d="M1487.445,132.809v24.403h-30.802v-24.403H1487.445z M1487.445,176.976v122.028h-30.802V176.976H1487.445z
			"/>
		<path fill="#FC7E00" d="M1547.291,132.809v166.195h-30.799V132.809H1547.291z"/>
		<path fill="#FC7E00" d="M1684.428,291.686c-18.672,4.887-36.905,7.318-54.736,7.318c-39.433,0-59.156-21.145-59.156-63.451
			c0-39.045,19.28-58.577,57.871-58.577c8.219,0,16.629,1.934,25.219,5.817v-49.984h30.803V291.686z M1653.625,208.83
			c-6.351-4.188-14.334-6.286-23.934-6.286c-19.129,0-28.717,10.731-28.717,32.197c0,25.494,9.975,38.244,29.877,38.244
			c8.053,0,15.646-1.135,22.773-3.369V208.83z"/>
		<path fill="#FC7E00" d="M1877.352,132.809v26.739h-47.653v139.456h-30.784V159.548h-47.652v-26.739H1877.352z"/>
		<path fill="#FC7E00" d="M1868.649,237.999c0-40.91,20.136-61.365,60.438-61.365c40.275,0,60.426,20.455,60.426,61.365
			c0,40.828-20.15,61.24-60.426,61.24C1888.949,299.239,1868.8,278.827,1868.649,237.999z M1929.088,275.772
			c19.751,0,29.627-12.75,29.627-38.244c0-24.877-9.876-37.304-29.627-37.304c-19.764,0-29.64,12.427-29.64,37.304
			C1899.448,263.022,1909.324,275.772,1929.088,275.772z"/>
		<path fill="#FC7E00" d="M2006.944,237.999c0-40.91,20.153-61.365,60.438-61.365c40.289,0,60.426,20.455,60.426,61.365
			c0,40.828-20.137,61.24-60.426,61.24C2027.248,299.239,2007.096,278.827,2006.944,237.999z M2067.383,275.772
			c19.768,0,29.627-12.75,29.627-38.244c0-24.877-9.859-37.304-29.627-37.304c-19.764,0-29.64,12.427-29.64,37.304
			C2037.743,263.022,2047.619,275.772,2067.383,275.772z"/>
		<path fill="#FC7E00" d="M2181.869,132.809v166.195h-30.799V132.809H2181.869z"/>
		<path fill="#FC7E00" d="M2210.915,293.202v-25.58c13.55,5.432,29.211,8.15,46.946,8.15c13.259,0,19.89-4.27,19.89-12.791
			c0-8.131-4.463-12.205-13.369-12.205h-22.086c-24.79,0-37.194-12.201-37.194-36.602c0-25.583,18.091-38.357,54.282-38.357
			c15.328,0,29.791,2.32,43.341,6.977v25.566c-13.55-5.43-28.273-8.136-44.157-8.136c-16.658,0-24.987,4.253-24.987,12.789
			c0,8.13,4.834,12.192,14.529,12.192h19.754c27.126,0,40.688,12.215,40.688,36.613c0,25.568-17.293,38.361-51.851,38.361
			C2239.74,300.18,2224.465,297.842,2210.915,293.202z"/>
	</g>
</g>
</svg>
